// Qsys_system.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module Qsys_system (
		input  wire        clk_clk,                     //                  clk.clk
		input  wire        pio_chaos_done_wire_export,  //  pio_chaos_done_wire.export
		output wire        pio_chaos_reset_wire_export, // pio_chaos_reset_wire.export
		output wire [31:0] pio_chaos_shift_wire_export, // pio_chaos_shift_wire.export
		output wire        pio_chaos_step_wire_export,  //  pio_chaos_step_wire.export
		input  wire [7:0]  pio_chaos_w_wire_export,     //     pio_chaos_w_wire.export
		input  wire [7:0]  pio_chaos_x_wire_export,     //     pio_chaos_x_wire.export
		input  wire [7:0]  pio_chaos_y_wire_export,     //     pio_chaos_y_wire.export
		input  wire [7:0]  pio_chaos_z_wire_export,     //     pio_chaos_z_wire.export
		input  wire        reset_reset_n,               //                reset.reset_n
		output wire        sdram_clk_clk,               //            sdram_clk.clk
		output wire [12:0] sdram_wire_addr,             //           sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,               //                     .ba
		output wire        sdram_wire_cas_n,            //                     .cas_n
		output wire        sdram_wire_cke,              //                     .cke
		output wire        sdram_wire_cs_n,             //                     .cs_n
		inout  wire [31:0] sdram_wire_dq,               //                     .dq
		output wire [3:0]  sdram_wire_dqm,              //                     .dqm
		output wire        sdram_wire_ras_n,            //                     .ras_n
		output wire        sdram_wire_we_n              //                     .we_n
	);

	wire         altpll_c0_clk;                                             // altpll:c0 -> [irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:altpll_c0_clk, nios2_gen2:clk, pio_chaos_done:clk, pio_chaos_reset:clk, pio_chaos_shift:clk, pio_chaos_step:clk, pio_chaos_w:clk, pio_chaos_x:clk, pio_chaos_y:clk, pio_chaos_z:clk, rst_controller_001:clk, sdram:clk, sysid:clock, timer:clk]
	wire  [31:0] nios2_gen2_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire         nios2_gen2_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire         nios2_gen2_data_master_debugaccess;                        // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire  [28:0] nios2_gen2_data_master_address;                            // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire   [3:0] nios2_gen2_data_master_byteenable;                         // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire         nios2_gen2_data_master_read;                               // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire         nios2_gen2_data_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_data_master_readdatavalid -> nios2_gen2:d_readdatavalid
	wire         nios2_gen2_data_master_write;                              // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire  [31:0] nios2_gen2_data_master_writedata;                          // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire  [31:0] nios2_gen2_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire         nios2_gen2_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire  [28:0] nios2_gen2_instruction_master_address;                     // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire         nios2_gen2_instruction_master_read;                        // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire         nios2_gen2_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;     // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;  // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_readdata;               // altpll:readdata -> mm_interconnect_0:altpll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_pll_slave_address;                // mm_interconnect_0:altpll_pll_slave_address -> altpll:address
	wire         mm_interconnect_0_altpll_pll_slave_read;                   // mm_interconnect_0:altpll_pll_slave_read -> altpll:read
	wire         mm_interconnect_0_altpll_pll_slave_write;                  // mm_interconnect_0:altpll_pll_slave_write -> altpll:write
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_writedata;              // mm_interconnect_0:altpll_pll_slave_writedata -> altpll:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_pio_chaos_step_s1_chipselect;            // mm_interconnect_0:pio_chaos_step_s1_chipselect -> pio_chaos_step:chipselect
	wire  [31:0] mm_interconnect_0_pio_chaos_step_s1_readdata;              // pio_chaos_step:readdata -> mm_interconnect_0:pio_chaos_step_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_chaos_step_s1_address;               // mm_interconnect_0:pio_chaos_step_s1_address -> pio_chaos_step:address
	wire         mm_interconnect_0_pio_chaos_step_s1_write;                 // mm_interconnect_0:pio_chaos_step_s1_write -> pio_chaos_step:write_n
	wire  [31:0] mm_interconnect_0_pio_chaos_step_s1_writedata;             // mm_interconnect_0:pio_chaos_step_s1_writedata -> pio_chaos_step:writedata
	wire         mm_interconnect_0_pio_chaos_reset_s1_chipselect;           // mm_interconnect_0:pio_chaos_reset_s1_chipselect -> pio_chaos_reset:chipselect
	wire  [31:0] mm_interconnect_0_pio_chaos_reset_s1_readdata;             // pio_chaos_reset:readdata -> mm_interconnect_0:pio_chaos_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_chaos_reset_s1_address;              // mm_interconnect_0:pio_chaos_reset_s1_address -> pio_chaos_reset:address
	wire         mm_interconnect_0_pio_chaos_reset_s1_write;                // mm_interconnect_0:pio_chaos_reset_s1_write -> pio_chaos_reset:write_n
	wire  [31:0] mm_interconnect_0_pio_chaos_reset_s1_writedata;            // mm_interconnect_0:pio_chaos_reset_s1_writedata -> pio_chaos_reset:writedata
	wire         mm_interconnect_0_pio_chaos_shift_s1_chipselect;           // mm_interconnect_0:pio_chaos_shift_s1_chipselect -> pio_chaos_shift:chipselect
	wire  [31:0] mm_interconnect_0_pio_chaos_shift_s1_readdata;             // pio_chaos_shift:readdata -> mm_interconnect_0:pio_chaos_shift_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_chaos_shift_s1_address;              // mm_interconnect_0:pio_chaos_shift_s1_address -> pio_chaos_shift:address
	wire         mm_interconnect_0_pio_chaos_shift_s1_write;                // mm_interconnect_0:pio_chaos_shift_s1_write -> pio_chaos_shift:write_n
	wire  [31:0] mm_interconnect_0_pio_chaos_shift_s1_writedata;            // mm_interconnect_0:pio_chaos_shift_s1_writedata -> pio_chaos_shift:writedata
	wire         mm_interconnect_0_pio_chaos_done_s1_chipselect;            // mm_interconnect_0:pio_chaos_done_s1_chipselect -> pio_chaos_done:chipselect
	wire  [31:0] mm_interconnect_0_pio_chaos_done_s1_readdata;              // pio_chaos_done:readdata -> mm_interconnect_0:pio_chaos_done_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_chaos_done_s1_address;               // mm_interconnect_0:pio_chaos_done_s1_address -> pio_chaos_done:address
	wire         mm_interconnect_0_pio_chaos_done_s1_write;                 // mm_interconnect_0:pio_chaos_done_s1_write -> pio_chaos_done:write_n
	wire  [31:0] mm_interconnect_0_pio_chaos_done_s1_writedata;             // mm_interconnect_0:pio_chaos_done_s1_writedata -> pio_chaos_done:writedata
	wire         mm_interconnect_0_pio_chaos_x_s1_chipselect;               // mm_interconnect_0:pio_chaos_x_s1_chipselect -> pio_chaos_x:chipselect
	wire  [31:0] mm_interconnect_0_pio_chaos_x_s1_readdata;                 // pio_chaos_x:readdata -> mm_interconnect_0:pio_chaos_x_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_chaos_x_s1_address;                  // mm_interconnect_0:pio_chaos_x_s1_address -> pio_chaos_x:address
	wire         mm_interconnect_0_pio_chaos_x_s1_write;                    // mm_interconnect_0:pio_chaos_x_s1_write -> pio_chaos_x:write_n
	wire  [31:0] mm_interconnect_0_pio_chaos_x_s1_writedata;                // mm_interconnect_0:pio_chaos_x_s1_writedata -> pio_chaos_x:writedata
	wire         mm_interconnect_0_pio_chaos_y_s1_chipselect;               // mm_interconnect_0:pio_chaos_y_s1_chipselect -> pio_chaos_y:chipselect
	wire  [31:0] mm_interconnect_0_pio_chaos_y_s1_readdata;                 // pio_chaos_y:readdata -> mm_interconnect_0:pio_chaos_y_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_chaos_y_s1_address;                  // mm_interconnect_0:pio_chaos_y_s1_address -> pio_chaos_y:address
	wire         mm_interconnect_0_pio_chaos_y_s1_write;                    // mm_interconnect_0:pio_chaos_y_s1_write -> pio_chaos_y:write_n
	wire  [31:0] mm_interconnect_0_pio_chaos_y_s1_writedata;                // mm_interconnect_0:pio_chaos_y_s1_writedata -> pio_chaos_y:writedata
	wire         mm_interconnect_0_pio_chaos_z_s1_chipselect;               // mm_interconnect_0:pio_chaos_z_s1_chipselect -> pio_chaos_z:chipselect
	wire  [31:0] mm_interconnect_0_pio_chaos_z_s1_readdata;                 // pio_chaos_z:readdata -> mm_interconnect_0:pio_chaos_z_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_chaos_z_s1_address;                  // mm_interconnect_0:pio_chaos_z_s1_address -> pio_chaos_z:address
	wire         mm_interconnect_0_pio_chaos_z_s1_write;                    // mm_interconnect_0:pio_chaos_z_s1_write -> pio_chaos_z:write_n
	wire  [31:0] mm_interconnect_0_pio_chaos_z_s1_writedata;                // mm_interconnect_0:pio_chaos_z_s1_writedata -> pio_chaos_z:writedata
	wire         mm_interconnect_0_pio_chaos_w_s1_chipselect;               // mm_interconnect_0:pio_chaos_w_s1_chipselect -> pio_chaos_w:chipselect
	wire  [31:0] mm_interconnect_0_pio_chaos_w_s1_readdata;                 // pio_chaos_w:readdata -> mm_interconnect_0:pio_chaos_w_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_chaos_w_s1_address;                  // mm_interconnect_0:pio_chaos_w_s1_address -> pio_chaos_w:address
	wire         mm_interconnect_0_pio_chaos_w_s1_write;                    // mm_interconnect_0:pio_chaos_w_s1_write -> pio_chaos_w:write_n
	wire  [31:0] mm_interconnect_0_pio_chaos_w_s1_writedata;                // mm_interconnect_0:pio_chaos_w_s1_writedata -> pio_chaos_w:writedata
	wire         irq_mapper_receiver0_irq;                                  // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [altpll:reset, mm_interconnect_0:altpll_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n, pio_chaos_done:reset_n, pio_chaos_reset:reset_n, pio_chaos_shift:reset_n, pio_chaos_step:reset_n, pio_chaos_w:reset_n, pio_chaos_x:reset_n, pio_chaos_y:reset_n, pio_chaos_z:reset_n, rst_translator:in_reset, sdram:reset_n, sysid:reset_n, timer:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [nios2_gen2:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_debug_reset_request_reset;                      // nios2_gen2:debug_reset_request -> rst_controller_001:reset_in1

	Qsys_system_altpll altpll (
		.clk       (clk_clk),                                      //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),               // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_pll_slave_writedata), //                      .writedata
		.c0        (altpll_c0_clk),                                //                    c0.clk
		.c1        (sdram_clk_clk),                                //                    c1.clk
		.areset    (),                                             //        areset_conduit.export
		.locked    (),                                             //        locked_conduit.export
		.phasedone ()                                              //     phasedone_conduit.export
	);

	Qsys_system_jtag_uart jtag_uart (
		.clk            (altpll_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	Qsys_system_nios2_gen2 nios2_gen2 (
		.clk                                 (altpll_c0_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	Qsys_system_pio_chaos_done pio_chaos_done (
		.clk        (altpll_c0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_chaos_done_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_chaos_done_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_chaos_done_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_chaos_done_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_chaos_done_s1_readdata),   //                    .readdata
		.in_port    (pio_chaos_done_wire_export)                      // external_connection.export
	);

	Qsys_system_pio_chaos_reset pio_chaos_reset (
		.clk        (altpll_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pio_chaos_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_chaos_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_chaos_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_chaos_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_chaos_reset_s1_readdata),   //                    .readdata
		.out_port   (pio_chaos_reset_wire_export)                      // external_connection.export
	);

	Qsys_system_pio_chaos_shift pio_chaos_shift (
		.clk        (altpll_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pio_chaos_shift_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_chaos_shift_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_chaos_shift_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_chaos_shift_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_chaos_shift_s1_readdata),   //                    .readdata
		.out_port   (pio_chaos_shift_wire_export)                      // external_connection.export
	);

	Qsys_system_pio_chaos_reset pio_chaos_step (
		.clk        (altpll_c0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_chaos_step_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_chaos_step_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_chaos_step_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_chaos_step_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_chaos_step_s1_readdata),   //                    .readdata
		.out_port   (pio_chaos_step_wire_export)                      // external_connection.export
	);

	Qsys_system_pio_chaos_w pio_chaos_w (
		.clk        (altpll_c0_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_chaos_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_chaos_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_chaos_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_chaos_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_chaos_w_s1_readdata),   //                    .readdata
		.in_port    (pio_chaos_w_wire_export)                      // external_connection.export
	);

	Qsys_system_pio_chaos_w pio_chaos_x (
		.clk        (altpll_c0_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_chaos_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_chaos_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_chaos_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_chaos_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_chaos_x_s1_readdata),   //                    .readdata
		.in_port    (pio_chaos_x_wire_export)                      // external_connection.export
	);

	Qsys_system_pio_chaos_w pio_chaos_y (
		.clk        (altpll_c0_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_chaos_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_chaos_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_chaos_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_chaos_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_chaos_y_s1_readdata),   //                    .readdata
		.in_port    (pio_chaos_y_wire_export)                      // external_connection.export
	);

	Qsys_system_pio_chaos_w pio_chaos_z (
		.clk        (altpll_c0_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_chaos_z_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_chaos_z_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_chaos_z_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_chaos_z_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_chaos_z_s1_readdata),   //                    .readdata
		.in_port    (pio_chaos_z_wire_export)                      // external_connection.export
	);

	Qsys_system_sdram sdram (
		.clk            (altpll_c0_clk),                            //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	Qsys_system_sysid sysid (
		.clock    (altpll_c0_clk),                                  //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	Qsys_system_timer timer (
		.clk        (altpll_c0_clk),                         //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	Qsys_system_mm_interconnect_0 mm_interconnect_0 (
		.altpll_c0_clk                                            (altpll_c0_clk),                                             //                                          altpll_c0.clk
		.clk_clk_clk                                              (clk_clk),                                                   //                                            clk_clk.clk
		.altpll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // altpll_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_gen2_reset_reset_bridge_in_reset_reset             (rst_controller_001_reset_out_reset),                        //             nios2_gen2_reset_reset_bridge_in_reset.reset
		.nios2_gen2_data_master_address                           (nios2_gen2_data_master_address),                            //                             nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                       (nios2_gen2_data_master_waitrequest),                        //                                                   .waitrequest
		.nios2_gen2_data_master_byteenable                        (nios2_gen2_data_master_byteenable),                         //                                                   .byteenable
		.nios2_gen2_data_master_read                              (nios2_gen2_data_master_read),                               //                                                   .read
		.nios2_gen2_data_master_readdata                          (nios2_gen2_data_master_readdata),                           //                                                   .readdata
		.nios2_gen2_data_master_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                      //                                                   .readdatavalid
		.nios2_gen2_data_master_write                             (nios2_gen2_data_master_write),                              //                                                   .write
		.nios2_gen2_data_master_writedata                         (nios2_gen2_data_master_writedata),                          //                                                   .writedata
		.nios2_gen2_data_master_debugaccess                       (nios2_gen2_data_master_debugaccess),                        //                                                   .debugaccess
		.nios2_gen2_instruction_master_address                    (nios2_gen2_instruction_master_address),                     //                      nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest                (nios2_gen2_instruction_master_waitrequest),                 //                                                   .waitrequest
		.nios2_gen2_instruction_master_read                       (nios2_gen2_instruction_master_read),                        //                                                   .read
		.nios2_gen2_instruction_master_readdata                   (nios2_gen2_instruction_master_readdata),                    //                                                   .readdata
		.nios2_gen2_instruction_master_readdatavalid              (nios2_gen2_instruction_master_readdatavalid),               //                                                   .readdatavalid
		.altpll_pll_slave_address                                 (mm_interconnect_0_altpll_pll_slave_address),                //                                   altpll_pll_slave.address
		.altpll_pll_slave_write                                   (mm_interconnect_0_altpll_pll_slave_write),                  //                                                   .write
		.altpll_pll_slave_read                                    (mm_interconnect_0_altpll_pll_slave_read),                   //                                                   .read
		.altpll_pll_slave_readdata                                (mm_interconnect_0_altpll_pll_slave_readdata),               //                                                   .readdata
		.altpll_pll_slave_writedata                               (mm_interconnect_0_altpll_pll_slave_writedata),              //                                                   .writedata
		.jtag_uart_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                   .write
		.jtag_uart_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                   .read
		.jtag_uart_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                   .chipselect
		.nios2_gen2_debug_mem_slave_address                       (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),      //                         nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                         (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),        //                                                   .write
		.nios2_gen2_debug_mem_slave_read                          (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),         //                                                   .read
		.nios2_gen2_debug_mem_slave_readdata                      (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),     //                                                   .readdata
		.nios2_gen2_debug_mem_slave_writedata                     (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),    //                                                   .writedata
		.nios2_gen2_debug_mem_slave_byteenable                    (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),   //                                                   .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest                   (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),  //                                                   .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess                   (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),  //                                                   .debugaccess
		.pio_chaos_done_s1_address                                (mm_interconnect_0_pio_chaos_done_s1_address),               //                                  pio_chaos_done_s1.address
		.pio_chaos_done_s1_write                                  (mm_interconnect_0_pio_chaos_done_s1_write),                 //                                                   .write
		.pio_chaos_done_s1_readdata                               (mm_interconnect_0_pio_chaos_done_s1_readdata),              //                                                   .readdata
		.pio_chaos_done_s1_writedata                              (mm_interconnect_0_pio_chaos_done_s1_writedata),             //                                                   .writedata
		.pio_chaos_done_s1_chipselect                             (mm_interconnect_0_pio_chaos_done_s1_chipselect),            //                                                   .chipselect
		.pio_chaos_reset_s1_address                               (mm_interconnect_0_pio_chaos_reset_s1_address),              //                                 pio_chaos_reset_s1.address
		.pio_chaos_reset_s1_write                                 (mm_interconnect_0_pio_chaos_reset_s1_write),                //                                                   .write
		.pio_chaos_reset_s1_readdata                              (mm_interconnect_0_pio_chaos_reset_s1_readdata),             //                                                   .readdata
		.pio_chaos_reset_s1_writedata                             (mm_interconnect_0_pio_chaos_reset_s1_writedata),            //                                                   .writedata
		.pio_chaos_reset_s1_chipselect                            (mm_interconnect_0_pio_chaos_reset_s1_chipselect),           //                                                   .chipselect
		.pio_chaos_shift_s1_address                               (mm_interconnect_0_pio_chaos_shift_s1_address),              //                                 pio_chaos_shift_s1.address
		.pio_chaos_shift_s1_write                                 (mm_interconnect_0_pio_chaos_shift_s1_write),                //                                                   .write
		.pio_chaos_shift_s1_readdata                              (mm_interconnect_0_pio_chaos_shift_s1_readdata),             //                                                   .readdata
		.pio_chaos_shift_s1_writedata                             (mm_interconnect_0_pio_chaos_shift_s1_writedata),            //                                                   .writedata
		.pio_chaos_shift_s1_chipselect                            (mm_interconnect_0_pio_chaos_shift_s1_chipselect),           //                                                   .chipselect
		.pio_chaos_step_s1_address                                (mm_interconnect_0_pio_chaos_step_s1_address),               //                                  pio_chaos_step_s1.address
		.pio_chaos_step_s1_write                                  (mm_interconnect_0_pio_chaos_step_s1_write),                 //                                                   .write
		.pio_chaos_step_s1_readdata                               (mm_interconnect_0_pio_chaos_step_s1_readdata),              //                                                   .readdata
		.pio_chaos_step_s1_writedata                              (mm_interconnect_0_pio_chaos_step_s1_writedata),             //                                                   .writedata
		.pio_chaos_step_s1_chipselect                             (mm_interconnect_0_pio_chaos_step_s1_chipselect),            //                                                   .chipselect
		.pio_chaos_w_s1_address                                   (mm_interconnect_0_pio_chaos_w_s1_address),                  //                                     pio_chaos_w_s1.address
		.pio_chaos_w_s1_write                                     (mm_interconnect_0_pio_chaos_w_s1_write),                    //                                                   .write
		.pio_chaos_w_s1_readdata                                  (mm_interconnect_0_pio_chaos_w_s1_readdata),                 //                                                   .readdata
		.pio_chaos_w_s1_writedata                                 (mm_interconnect_0_pio_chaos_w_s1_writedata),                //                                                   .writedata
		.pio_chaos_w_s1_chipselect                                (mm_interconnect_0_pio_chaos_w_s1_chipselect),               //                                                   .chipselect
		.pio_chaos_x_s1_address                                   (mm_interconnect_0_pio_chaos_x_s1_address),                  //                                     pio_chaos_x_s1.address
		.pio_chaos_x_s1_write                                     (mm_interconnect_0_pio_chaos_x_s1_write),                    //                                                   .write
		.pio_chaos_x_s1_readdata                                  (mm_interconnect_0_pio_chaos_x_s1_readdata),                 //                                                   .readdata
		.pio_chaos_x_s1_writedata                                 (mm_interconnect_0_pio_chaos_x_s1_writedata),                //                                                   .writedata
		.pio_chaos_x_s1_chipselect                                (mm_interconnect_0_pio_chaos_x_s1_chipselect),               //                                                   .chipselect
		.pio_chaos_y_s1_address                                   (mm_interconnect_0_pio_chaos_y_s1_address),                  //                                     pio_chaos_y_s1.address
		.pio_chaos_y_s1_write                                     (mm_interconnect_0_pio_chaos_y_s1_write),                    //                                                   .write
		.pio_chaos_y_s1_readdata                                  (mm_interconnect_0_pio_chaos_y_s1_readdata),                 //                                                   .readdata
		.pio_chaos_y_s1_writedata                                 (mm_interconnect_0_pio_chaos_y_s1_writedata),                //                                                   .writedata
		.pio_chaos_y_s1_chipselect                                (mm_interconnect_0_pio_chaos_y_s1_chipselect),               //                                                   .chipselect
		.pio_chaos_z_s1_address                                   (mm_interconnect_0_pio_chaos_z_s1_address),                  //                                     pio_chaos_z_s1.address
		.pio_chaos_z_s1_write                                     (mm_interconnect_0_pio_chaos_z_s1_write),                    //                                                   .write
		.pio_chaos_z_s1_readdata                                  (mm_interconnect_0_pio_chaos_z_s1_readdata),                 //                                                   .readdata
		.pio_chaos_z_s1_writedata                                 (mm_interconnect_0_pio_chaos_z_s1_writedata),                //                                                   .writedata
		.pio_chaos_z_s1_chipselect                                (mm_interconnect_0_pio_chaos_z_s1_chipselect),               //                                                   .chipselect
		.sdram_s1_address                                         (mm_interconnect_0_sdram_s1_address),                        //                                           sdram_s1.address
		.sdram_s1_write                                           (mm_interconnect_0_sdram_s1_write),                          //                                                   .write
		.sdram_s1_read                                            (mm_interconnect_0_sdram_s1_read),                           //                                                   .read
		.sdram_s1_readdata                                        (mm_interconnect_0_sdram_s1_readdata),                       //                                                   .readdata
		.sdram_s1_writedata                                       (mm_interconnect_0_sdram_s1_writedata),                      //                                                   .writedata
		.sdram_s1_byteenable                                      (mm_interconnect_0_sdram_s1_byteenable),                     //                                                   .byteenable
		.sdram_s1_readdatavalid                                   (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                                   .readdatavalid
		.sdram_s1_waitrequest                                     (mm_interconnect_0_sdram_s1_waitrequest),                    //                                                   .waitrequest
		.sdram_s1_chipselect                                      (mm_interconnect_0_sdram_s1_chipselect),                     //                                                   .chipselect
		.sysid_control_slave_address                              (mm_interconnect_0_sysid_control_slave_address),             //                                sysid_control_slave.address
		.sysid_control_slave_readdata                             (mm_interconnect_0_sysid_control_slave_readdata),            //                                                   .readdata
		.timer_s1_address                                         (mm_interconnect_0_timer_s1_address),                        //                                           timer_s1.address
		.timer_s1_write                                           (mm_interconnect_0_timer_s1_write),                          //                                                   .write
		.timer_s1_readdata                                        (mm_interconnect_0_timer_s1_readdata),                       //                                                   .readdata
		.timer_s1_writedata                                       (mm_interconnect_0_timer_s1_writedata),                      //                                                   .writedata
		.timer_s1_chipselect                                      (mm_interconnect_0_timer_s1_chipselect)                      //                                                   .chipselect
	);

	Qsys_system_irq_mapper irq_mapper (
		.clk           (altpll_c0_clk),                      //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_gen2_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset),   // reset_in1.reset
		.clk            (altpll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
