// Qsys_system.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module Qsys_system (
		input  wire        chaos_code_done_wire_export,  //  chaos_code_done_wire.export
		output wire        chaos_code_reset_wire_export, // chaos_code_reset_wire.export
		output wire [31:0] chaos_code_shift_wire_export, // chaos_code_shift_wire.export
		output wire        chaos_code_step_wire_export,  //  chaos_code_step_wire.export
		input  wire [7:0]  chaos_code_w_wire_export,     //     chaos_code_w_wire.export
		input  wire [7:0]  chaos_code_x_wire_export,     //     chaos_code_x_wire.export
		input  wire [7:0]  chaos_code_y_wire_export,     //     chaos_code_y_wire.export
		input  wire [7:0]  chaos_code_z_wire_export,     //     chaos_code_z_wire.export
		input  wire        clk_clk,                      //                   clk.clk
		input  wire [1:0]  pio_key_wire_export,          //          pio_key_wire.export
		output wire [3:0]  pio_led_wire_export,          //          pio_led_wire.export
		output wire        pio_wifi_reset_wire_export,   //   pio_wifi_reset_wire.export
		inout  wire [15:0] pixel_buffer_wire_DQ,         //     pixel_buffer_wire.DQ
		output wire [19:0] pixel_buffer_wire_ADDR,       //                      .ADDR
		output wire        pixel_buffer_wire_LB_N,       //                      .LB_N
		output wire        pixel_buffer_wire_UB_N,       //                      .UB_N
		output wire        pixel_buffer_wire_CE_N,       //                      .CE_N
		output wire        pixel_buffer_wire_OE_N,       //                      .OE_N
		output wire        pixel_buffer_wire_WE_N,       //                      .WE_N
		input  wire        reset_reset_n,                //                 reset.reset_n
		inout  wire        sd_card_wire_b_SD_cmd,        //          sd_card_wire.b_SD_cmd
		inout  wire        sd_card_wire_b_SD_dat,        //                      .b_SD_dat
		inout  wire        sd_card_wire_b_SD_dat3,       //                      .b_SD_dat3
		output wire        sd_card_wire_o_SD_clock,      //                      .o_SD_clock
		output wire        sdram_clk_clk,                //             sdram_clk.clk
		output wire [12:0] sdram_wire_addr,              //            sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                //                      .ba
		output wire        sdram_wire_cas_n,             //                      .cas_n
		output wire        sdram_wire_cke,               //                      .cke
		output wire        sdram_wire_cs_n,              //                      .cs_n
		inout  wire [31:0] sdram_wire_dq,                //                      .dq
		output wire [3:0]  sdram_wire_dqm,               //                      .dqm
		output wire        sdram_wire_ras_n,             //                      .ras_n
		output wire        sdram_wire_we_n,              //                      .we_n
		output wire        vga_controller_wire_CLK,      //   vga_controller_wire.CLK
		output wire        vga_controller_wire_HS,       //                      .HS
		output wire        vga_controller_wire_VS,       //                      .VS
		output wire        vga_controller_wire_BLANK,    //                      .BLANK
		output wire        vga_controller_wire_SYNC,     //                      .SYNC
		output wire [7:0]  vga_controller_wire_R,        //                      .R
		output wire [7:0]  vga_controller_wire_G,        //                      .G
		output wire [7:0]  vga_controller_wire_B,        //                      .B
		input  wire        wifi_uart_wire_rxd,           //        wifi_uart_wire.rxd
		output wire        wifi_uart_wire_txd,           //                      .txd
		input  wire        wifi_uart_wire_cts_n,         //                      .cts_n
		output wire        wifi_uart_wire_rts_n          //                      .rts_n
	);

	wire         dual_clock_buffer_avalon_dc_buffer_source_valid;                    // dual_clock_buffer:stream_out_valid -> vga_controller:valid
	wire  [29:0] dual_clock_buffer_avalon_dc_buffer_source_data;                     // dual_clock_buffer:stream_out_data -> vga_controller:data
	wire         dual_clock_buffer_avalon_dc_buffer_source_ready;                    // vga_controller:ready -> dual_clock_buffer:stream_out_ready
	wire         dual_clock_buffer_avalon_dc_buffer_source_startofpacket;            // dual_clock_buffer:stream_out_startofpacket -> vga_controller:startofpacket
	wire         dual_clock_buffer_avalon_dc_buffer_source_endofpacket;              // dual_clock_buffer:stream_out_endofpacket -> vga_controller:endofpacket
	wire         pixel_buffer_dma_avalon_pixel_source_valid;                         // pixel_buffer_dma:stream_valid -> video_rgb_resampler_0:stream_in_valid
	wire  [23:0] pixel_buffer_dma_avalon_pixel_source_data;                          // pixel_buffer_dma:stream_data -> video_rgb_resampler_0:stream_in_data
	wire         pixel_buffer_dma_avalon_pixel_source_ready;                         // video_rgb_resampler_0:stream_in_ready -> pixel_buffer_dma:stream_ready
	wire         pixel_buffer_dma_avalon_pixel_source_startofpacket;                 // pixel_buffer_dma:stream_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire         pixel_buffer_dma_avalon_pixel_source_endofpacket;                   // pixel_buffer_dma:stream_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_valid;                      // video_rgb_resampler_0:stream_out_valid -> dual_clock_buffer:stream_in_valid
	wire  [29:0] video_rgb_resampler_0_avalon_rgb_source_data;                       // video_rgb_resampler_0:stream_out_data -> dual_clock_buffer:stream_in_data
	wire         video_rgb_resampler_0_avalon_rgb_source_ready;                      // dual_clock_buffer:stream_in_ready -> video_rgb_resampler_0:stream_out_ready
	wire         video_rgb_resampler_0_avalon_rgb_source_startofpacket;              // video_rgb_resampler_0:stream_out_startofpacket -> dual_clock_buffer:stream_in_startofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_endofpacket;                // video_rgb_resampler_0:stream_out_endofpacket -> dual_clock_buffer:stream_in_endofpacket
	wire         altpll_c0_clk;                                                      // altpll:c0 -> [chaos_code_done:clk, chaos_code_reset:clk, chaos_code_shift:clk, chaos_code_step:clk, chaos_code_w:clk, chaos_code_x:clk, chaos_code_y:clk, chaos_code_z:clk, dual_clock_buffer:clk_stream_in, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:altpll_c0_clk, nios2_gen2:clk, pio_key:clk, pio_led:clk, pio_wifi_reset:clk, pixel_buffer:clk, pixel_buffer_dma:clk, rst_controller_001:clk, sd_card:i_clock, sdram:clk, sysid:clock, timer:clk, video_rgb_resampler_0:clk, wifi_uart:clk]
	wire         altpll_c2_clk;                                                      // altpll:c2 -> [dual_clock_buffer:clk_stream_out, rst_controller_002:clk, vga_controller:clk]
	wire         pixel_buffer_dma_avalon_pixel_dma_master_waitrequest;               // mm_interconnect_0:pixel_buffer_dma_avalon_pixel_dma_master_waitrequest -> pixel_buffer_dma:master_waitrequest
	wire  [31:0] pixel_buffer_dma_avalon_pixel_dma_master_readdata;                  // mm_interconnect_0:pixel_buffer_dma_avalon_pixel_dma_master_readdata -> pixel_buffer_dma:master_readdata
	wire  [31:0] pixel_buffer_dma_avalon_pixel_dma_master_address;                   // pixel_buffer_dma:master_address -> mm_interconnect_0:pixel_buffer_dma_avalon_pixel_dma_master_address
	wire         pixel_buffer_dma_avalon_pixel_dma_master_read;                      // pixel_buffer_dma:master_read -> mm_interconnect_0:pixel_buffer_dma_avalon_pixel_dma_master_read
	wire         pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid;             // mm_interconnect_0:pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid -> pixel_buffer_dma:master_readdatavalid
	wire         pixel_buffer_dma_avalon_pixel_dma_master_lock;                      // pixel_buffer_dma:master_arbiterlock -> mm_interconnect_0:pixel_buffer_dma_avalon_pixel_dma_master_lock
	wire  [31:0] nios2_gen2_data_master_readdata;                                    // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire         nios2_gen2_data_master_waitrequest;                                 // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire         nios2_gen2_data_master_debugaccess;                                 // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire  [28:0] nios2_gen2_data_master_address;                                     // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire   [3:0] nios2_gen2_data_master_byteenable;                                  // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire         nios2_gen2_data_master_read;                                        // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire         nios2_gen2_data_master_readdatavalid;                               // mm_interconnect_0:nios2_gen2_data_master_readdatavalid -> nios2_gen2:d_readdatavalid
	wire         nios2_gen2_data_master_write;                                       // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire  [31:0] nios2_gen2_data_master_writedata;                                   // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire  [31:0] nios2_gen2_instruction_master_readdata;                             // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire         nios2_gen2_instruction_master_waitrequest;                          // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire  [28:0] nios2_gen2_instruction_master_address;                              // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire         nios2_gen2_instruction_master_read;                                 // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire         nios2_gen2_instruction_master_readdatavalid;                        // mm_interconnect_0:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire  [15:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdata;          // pixel_buffer:readdata -> mm_interconnect_0:pixel_buffer_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_address;           // mm_interconnect_0:pixel_buffer_avalon_sram_slave_address -> pixel_buffer:address
	wire         mm_interconnect_0_pixel_buffer_avalon_sram_slave_read;              // mm_interconnect_0:pixel_buffer_avalon_sram_slave_read -> pixel_buffer:read
	wire   [1:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_byteenable;        // mm_interconnect_0:pixel_buffer_avalon_sram_slave_byteenable -> pixel_buffer:byteenable
	wire         mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdatavalid;     // pixel_buffer:readdatavalid -> mm_interconnect_0:pixel_buffer_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_pixel_buffer_avalon_sram_slave_write;             // mm_interconnect_0:pixel_buffer_avalon_sram_slave_write -> pixel_buffer:write
	wire  [15:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_writedata;         // mm_interconnect_0:pixel_buffer_avalon_sram_slave_writedata -> pixel_buffer:writedata
	wire  [31:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata;   // pixel_buffer_dma:slave_readdata -> mm_interconnect_0:pixel_buffer_dma_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address;    // mm_interconnect_0:pixel_buffer_dma_avalon_control_slave_address -> pixel_buffer_dma:slave_address
	wire         mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read;       // mm_interconnect_0:pixel_buffer_dma_avalon_control_slave_read -> pixel_buffer_dma:slave_read
	wire   [3:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable; // mm_interconnect_0:pixel_buffer_dma_avalon_control_slave_byteenable -> pixel_buffer_dma:slave_byteenable
	wire         mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write;      // mm_interconnect_0:pixel_buffer_dma_avalon_control_slave_write -> pixel_buffer_dma:slave_write
	wire  [31:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata;  // mm_interconnect_0:pixel_buffer_dma_avalon_control_slave_writedata -> pixel_buffer_dma:slave_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;             // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;          // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect;           // mm_interconnect_0:sd_card_avalon_sdcard_slave_chipselect -> sd_card:i_avalon_chip_select
	wire  [31:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata;             // sd_card:o_avalon_readdata -> mm_interconnect_0:sd_card_avalon_sdcard_slave_readdata
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest;          // sd_card:o_avalon_waitrequest -> mm_interconnect_0:sd_card_avalon_sdcard_slave_waitrequest
	wire   [7:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_address;              // mm_interconnect_0:sd_card_avalon_sdcard_slave_address -> sd_card:i_avalon_address
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_read;                 // mm_interconnect_0:sd_card_avalon_sdcard_slave_read -> sd_card:i_avalon_read
	wire   [3:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable;           // mm_interconnect_0:sd_card_avalon_sdcard_slave_byteenable -> sd_card:i_avalon_byteenable
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_write;                // mm_interconnect_0:sd_card_avalon_sdcard_slave_write -> sd_card:i_avalon_write
	wire  [31:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata;            // mm_interconnect_0:sd_card_avalon_sdcard_slave_writedata -> sd_card:i_avalon_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                     // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                      // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;              // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;           // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;           // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;               // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_read;                  // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;            // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_write;                 // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;             // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_readdata;                        // altpll:readdata -> mm_interconnect_0:altpll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_pll_slave_address;                         // mm_interconnect_0:altpll_pll_slave_address -> altpll:address
	wire         mm_interconnect_0_altpll_pll_slave_read;                            // mm_interconnect_0:altpll_pll_slave_read -> altpll:read
	wire         mm_interconnect_0_altpll_pll_slave_write;                           // mm_interconnect_0:altpll_pll_slave_write -> altpll:write
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_writedata;                       // mm_interconnect_0:altpll_pll_slave_writedata -> altpll:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                              // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                                // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                             // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                 // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                    // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                              // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                           // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                   // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                               // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_s1_chipselect;                              // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                                // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                 // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                   // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                               // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_wifi_uart_s1_chipselect;                          // mm_interconnect_0:wifi_uart_s1_chipselect -> wifi_uart:chipselect
	wire  [15:0] mm_interconnect_0_wifi_uart_s1_readdata;                            // wifi_uart:readdata -> mm_interconnect_0:wifi_uart_s1_readdata
	wire   [2:0] mm_interconnect_0_wifi_uart_s1_address;                             // mm_interconnect_0:wifi_uart_s1_address -> wifi_uart:address
	wire         mm_interconnect_0_wifi_uart_s1_read;                                // mm_interconnect_0:wifi_uart_s1_read -> wifi_uart:read_n
	wire         mm_interconnect_0_wifi_uart_s1_begintransfer;                       // mm_interconnect_0:wifi_uart_s1_begintransfer -> wifi_uart:begintransfer
	wire         mm_interconnect_0_wifi_uart_s1_write;                               // mm_interconnect_0:wifi_uart_s1_write -> wifi_uart:write_n
	wire  [15:0] mm_interconnect_0_wifi_uart_s1_writedata;                           // mm_interconnect_0:wifi_uart_s1_writedata -> wifi_uart:writedata
	wire         mm_interconnect_0_pio_wifi_reset_s1_chipselect;                     // mm_interconnect_0:pio_wifi_reset_s1_chipselect -> pio_wifi_reset:chipselect
	wire  [31:0] mm_interconnect_0_pio_wifi_reset_s1_readdata;                       // pio_wifi_reset:readdata -> mm_interconnect_0:pio_wifi_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_wifi_reset_s1_address;                        // mm_interconnect_0:pio_wifi_reset_s1_address -> pio_wifi_reset:address
	wire         mm_interconnect_0_pio_wifi_reset_s1_write;                          // mm_interconnect_0:pio_wifi_reset_s1_write -> pio_wifi_reset:write_n
	wire  [31:0] mm_interconnect_0_pio_wifi_reset_s1_writedata;                      // mm_interconnect_0:pio_wifi_reset_s1_writedata -> pio_wifi_reset:writedata
	wire         mm_interconnect_0_pio_led_s1_chipselect;                            // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                              // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                               // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_write;                                 // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                             // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire         mm_interconnect_0_pio_key_s1_chipselect;                            // mm_interconnect_0:pio_key_s1_chipselect -> pio_key:chipselect
	wire  [31:0] mm_interconnect_0_pio_key_s1_readdata;                              // pio_key:readdata -> mm_interconnect_0:pio_key_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_key_s1_address;                               // mm_interconnect_0:pio_key_s1_address -> pio_key:address
	wire         mm_interconnect_0_pio_key_s1_write;                                 // mm_interconnect_0:pio_key_s1_write -> pio_key:write_n
	wire  [31:0] mm_interconnect_0_pio_key_s1_writedata;                             // mm_interconnect_0:pio_key_s1_writedata -> pio_key:writedata
	wire         mm_interconnect_0_chaos_code_step_s1_chipselect;                    // mm_interconnect_0:chaos_code_step_s1_chipselect -> chaos_code_step:chipselect
	wire  [31:0] mm_interconnect_0_chaos_code_step_s1_readdata;                      // chaos_code_step:readdata -> mm_interconnect_0:chaos_code_step_s1_readdata
	wire   [1:0] mm_interconnect_0_chaos_code_step_s1_address;                       // mm_interconnect_0:chaos_code_step_s1_address -> chaos_code_step:address
	wire         mm_interconnect_0_chaos_code_step_s1_write;                         // mm_interconnect_0:chaos_code_step_s1_write -> chaos_code_step:write_n
	wire  [31:0] mm_interconnect_0_chaos_code_step_s1_writedata;                     // mm_interconnect_0:chaos_code_step_s1_writedata -> chaos_code_step:writedata
	wire         mm_interconnect_0_chaos_code_reset_s1_chipselect;                   // mm_interconnect_0:chaos_code_reset_s1_chipselect -> chaos_code_reset:chipselect
	wire  [31:0] mm_interconnect_0_chaos_code_reset_s1_readdata;                     // chaos_code_reset:readdata -> mm_interconnect_0:chaos_code_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_chaos_code_reset_s1_address;                      // mm_interconnect_0:chaos_code_reset_s1_address -> chaos_code_reset:address
	wire         mm_interconnect_0_chaos_code_reset_s1_write;                        // mm_interconnect_0:chaos_code_reset_s1_write -> chaos_code_reset:write_n
	wire  [31:0] mm_interconnect_0_chaos_code_reset_s1_writedata;                    // mm_interconnect_0:chaos_code_reset_s1_writedata -> chaos_code_reset:writedata
	wire         mm_interconnect_0_chaos_code_shift_s1_chipselect;                   // mm_interconnect_0:chaos_code_shift_s1_chipselect -> chaos_code_shift:chipselect
	wire  [31:0] mm_interconnect_0_chaos_code_shift_s1_readdata;                     // chaos_code_shift:readdata -> mm_interconnect_0:chaos_code_shift_s1_readdata
	wire   [1:0] mm_interconnect_0_chaos_code_shift_s1_address;                      // mm_interconnect_0:chaos_code_shift_s1_address -> chaos_code_shift:address
	wire         mm_interconnect_0_chaos_code_shift_s1_write;                        // mm_interconnect_0:chaos_code_shift_s1_write -> chaos_code_shift:write_n
	wire  [31:0] mm_interconnect_0_chaos_code_shift_s1_writedata;                    // mm_interconnect_0:chaos_code_shift_s1_writedata -> chaos_code_shift:writedata
	wire         mm_interconnect_0_chaos_code_done_s1_chipselect;                    // mm_interconnect_0:chaos_code_done_s1_chipselect -> chaos_code_done:chipselect
	wire  [31:0] mm_interconnect_0_chaos_code_done_s1_readdata;                      // chaos_code_done:readdata -> mm_interconnect_0:chaos_code_done_s1_readdata
	wire   [1:0] mm_interconnect_0_chaos_code_done_s1_address;                       // mm_interconnect_0:chaos_code_done_s1_address -> chaos_code_done:address
	wire         mm_interconnect_0_chaos_code_done_s1_write;                         // mm_interconnect_0:chaos_code_done_s1_write -> chaos_code_done:write_n
	wire  [31:0] mm_interconnect_0_chaos_code_done_s1_writedata;                     // mm_interconnect_0:chaos_code_done_s1_writedata -> chaos_code_done:writedata
	wire         mm_interconnect_0_chaos_code_x_s1_chipselect;                       // mm_interconnect_0:chaos_code_x_s1_chipselect -> chaos_code_x:chipselect
	wire  [31:0] mm_interconnect_0_chaos_code_x_s1_readdata;                         // chaos_code_x:readdata -> mm_interconnect_0:chaos_code_x_s1_readdata
	wire   [1:0] mm_interconnect_0_chaos_code_x_s1_address;                          // mm_interconnect_0:chaos_code_x_s1_address -> chaos_code_x:address
	wire         mm_interconnect_0_chaos_code_x_s1_write;                            // mm_interconnect_0:chaos_code_x_s1_write -> chaos_code_x:write_n
	wire  [31:0] mm_interconnect_0_chaos_code_x_s1_writedata;                        // mm_interconnect_0:chaos_code_x_s1_writedata -> chaos_code_x:writedata
	wire         mm_interconnect_0_chaos_code_y_s1_chipselect;                       // mm_interconnect_0:chaos_code_y_s1_chipselect -> chaos_code_y:chipselect
	wire  [31:0] mm_interconnect_0_chaos_code_y_s1_readdata;                         // chaos_code_y:readdata -> mm_interconnect_0:chaos_code_y_s1_readdata
	wire   [1:0] mm_interconnect_0_chaos_code_y_s1_address;                          // mm_interconnect_0:chaos_code_y_s1_address -> chaos_code_y:address
	wire         mm_interconnect_0_chaos_code_y_s1_write;                            // mm_interconnect_0:chaos_code_y_s1_write -> chaos_code_y:write_n
	wire  [31:0] mm_interconnect_0_chaos_code_y_s1_writedata;                        // mm_interconnect_0:chaos_code_y_s1_writedata -> chaos_code_y:writedata
	wire         mm_interconnect_0_chaos_code_z_s1_chipselect;                       // mm_interconnect_0:chaos_code_z_s1_chipselect -> chaos_code_z:chipselect
	wire  [31:0] mm_interconnect_0_chaos_code_z_s1_readdata;                         // chaos_code_z:readdata -> mm_interconnect_0:chaos_code_z_s1_readdata
	wire   [1:0] mm_interconnect_0_chaos_code_z_s1_address;                          // mm_interconnect_0:chaos_code_z_s1_address -> chaos_code_z:address
	wire         mm_interconnect_0_chaos_code_z_s1_write;                            // mm_interconnect_0:chaos_code_z_s1_write -> chaos_code_z:write_n
	wire  [31:0] mm_interconnect_0_chaos_code_z_s1_writedata;                        // mm_interconnect_0:chaos_code_z_s1_writedata -> chaos_code_z:writedata
	wire         mm_interconnect_0_chaos_code_w_s1_chipselect;                       // mm_interconnect_0:chaos_code_w_s1_chipselect -> chaos_code_w:chipselect
	wire  [31:0] mm_interconnect_0_chaos_code_w_s1_readdata;                         // chaos_code_w:readdata -> mm_interconnect_0:chaos_code_w_s1_readdata
	wire   [1:0] mm_interconnect_0_chaos_code_w_s1_address;                          // mm_interconnect_0:chaos_code_w_s1_address -> chaos_code_w:address
	wire         mm_interconnect_0_chaos_code_w_s1_write;                            // mm_interconnect_0:chaos_code_w_s1_write -> chaos_code_w:write_n
	wire  [31:0] mm_interconnect_0_chaos_code_w_s1_writedata;                        // mm_interconnect_0:chaos_code_w_s1_writedata -> chaos_code_w:writedata
	wire         irq_mapper_receiver0_irq;                                           // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                           // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                           // wifi_uart:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                           // pio_key:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_irq_irq;                                                 // irq_mapper:sender_irq -> nios2_gen2:irq
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [altpll:reset, mm_interconnect_0:altpll_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> [chaos_code_done:reset_n, chaos_code_reset:reset_n, chaos_code_shift:reset_n, chaos_code_step:reset_n, chaos_code_w:reset_n, chaos_code_x:reset_n, chaos_code_y:reset_n, chaos_code_z:reset_n, dual_clock_buffer:reset_stream_in, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:pixel_buffer_dma_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n, pio_key:reset_n, pio_led:reset_n, pio_wifi_reset:reset_n, pixel_buffer:reset, pixel_buffer_dma:reset, rst_translator:in_reset, sd_card:i_reset_n, sdram:reset_n, sysid:reset_n, timer:reset_n, video_rgb_resampler_0:reset, wifi_uart:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                             // rst_controller_001:reset_req -> [nios2_gen2:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_debug_reset_request_reset;                               // nios2_gen2:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                                 // rst_controller_002:reset_out -> [dual_clock_buffer:reset_stream_out, vga_controller:reset]

	Qsys_system_altpll altpll (
		.clk       (clk_clk),                                      //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),               // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_pll_slave_writedata), //                      .writedata
		.c0        (altpll_c0_clk),                                //                    c0.clk
		.c1        (sdram_clk_clk),                                //                    c1.clk
		.c2        (altpll_c2_clk),                                //                    c2.clk
		.areset    (),                                             //        areset_conduit.export
		.locked    (),                                             //        locked_conduit.export
		.phasedone ()                                              //     phasedone_conduit.export
	);

	Qsys_system_chaos_code_done chaos_code_done (
		.clk        (altpll_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_chaos_code_done_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chaos_code_done_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chaos_code_done_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chaos_code_done_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chaos_code_done_s1_readdata),   //                    .readdata
		.in_port    (chaos_code_done_wire_export)                      // external_connection.export
	);

	Qsys_system_chaos_code_reset chaos_code_reset (
		.clk        (altpll_c0_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chaos_code_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chaos_code_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chaos_code_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chaos_code_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chaos_code_reset_s1_readdata),   //                    .readdata
		.out_port   (chaos_code_reset_wire_export)                      // external_connection.export
	);

	Qsys_system_chaos_code_shift chaos_code_shift (
		.clk        (altpll_c0_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chaos_code_shift_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chaos_code_shift_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chaos_code_shift_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chaos_code_shift_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chaos_code_shift_s1_readdata),   //                    .readdata
		.out_port   (chaos_code_shift_wire_export)                      // external_connection.export
	);

	Qsys_system_chaos_code_reset chaos_code_step (
		.clk        (altpll_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_chaos_code_step_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chaos_code_step_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chaos_code_step_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chaos_code_step_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chaos_code_step_s1_readdata),   //                    .readdata
		.out_port   (chaos_code_step_wire_export)                      // external_connection.export
	);

	Qsys_system_chaos_code_w chaos_code_w (
		.clk        (altpll_c0_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_chaos_code_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chaos_code_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chaos_code_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chaos_code_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chaos_code_w_s1_readdata),   //                    .readdata
		.in_port    (chaos_code_w_wire_export)                      // external_connection.export
	);

	Qsys_system_chaos_code_w chaos_code_x (
		.clk        (altpll_c0_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_chaos_code_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chaos_code_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chaos_code_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chaos_code_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chaos_code_x_s1_readdata),   //                    .readdata
		.in_port    (chaos_code_x_wire_export)                      // external_connection.export
	);

	Qsys_system_chaos_code_w chaos_code_y (
		.clk        (altpll_c0_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_chaos_code_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chaos_code_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chaos_code_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chaos_code_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chaos_code_y_s1_readdata),   //                    .readdata
		.in_port    (chaos_code_y_wire_export)                      // external_connection.export
	);

	Qsys_system_chaos_code_w chaos_code_z (
		.clk        (altpll_c0_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_chaos_code_z_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chaos_code_z_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chaos_code_z_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chaos_code_z_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chaos_code_z_s1_readdata),   //                    .readdata
		.in_port    (chaos_code_z_wire_export)                      // external_connection.export
	);

	Qsys_system_dual_clock_buffer dual_clock_buffer (
		.clk_stream_in            (altpll_c0_clk),                                           //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_001_reset_out_reset),                      //         reset_stream_in.reset
		.clk_stream_out           (altpll_c2_clk),                                           //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                      //        reset_stream_out.reset
		.stream_in_ready          (video_rgb_resampler_0_avalon_rgb_source_ready),           //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (video_rgb_resampler_0_avalon_rgb_source_startofpacket),   //                        .startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_0_avalon_rgb_source_endofpacket),     //                        .endofpacket
		.stream_in_valid          (video_rgb_resampler_0_avalon_rgb_source_valid),           //                        .valid
		.stream_in_data           (video_rgb_resampler_0_avalon_rgb_source_data),            //                        .data
		.stream_out_ready         (dual_clock_buffer_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (dual_clock_buffer_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (dual_clock_buffer_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (dual_clock_buffer_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (dual_clock_buffer_avalon_dc_buffer_source_data)           //                        .data
	);

	Qsys_system_jtag_uart jtag_uart (
		.clk            (altpll_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	Qsys_system_nios2_gen2 nios2_gen2 (
		.clk                                 (altpll_c0_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	Qsys_system_pio_key pio_key (
		.clk        (altpll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_pio_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_key_s1_readdata),   //                    .readdata
		.in_port    (pio_key_wire_export),                     // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                 //                 irq.irq
	);

	Qsys_system_pio_led pio_led (
		.clk        (altpll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_wire_export)                      // external_connection.export
	);

	Qsys_system_pio_wifi_reset pio_wifi_reset (
		.clk        (altpll_c0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_wifi_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_wifi_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_wifi_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_wifi_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_wifi_reset_s1_readdata),   //                    .readdata
		.out_port   (pio_wifi_reset_wire_export)                      // external_connection.export
	);

	Qsys_system_pixel_buffer pixel_buffer (
		.clk           (altpll_c0_clk),                                                  //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),                             //              reset.reset
		.SRAM_DQ       (pixel_buffer_wire_DQ),                                           // external_interface.export
		.SRAM_ADDR     (pixel_buffer_wire_ADDR),                                         //                   .export
		.SRAM_LB_N     (pixel_buffer_wire_LB_N),                                         //                   .export
		.SRAM_UB_N     (pixel_buffer_wire_UB_N),                                         //                   .export
		.SRAM_CE_N     (pixel_buffer_wire_CE_N),                                         //                   .export
		.SRAM_OE_N     (pixel_buffer_wire_OE_N),                                         //                   .export
		.SRAM_WE_N     (pixel_buffer_wire_WE_N),                                         //                   .export
		.address       (mm_interconnect_0_pixel_buffer_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_pixel_buffer_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_pixel_buffer_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_pixel_buffer_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_pixel_buffer_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	Qsys_system_pixel_buffer_dma pixel_buffer_dma (
		.clk                  (altpll_c0_clk),                                                      //                     clk.clk
		.reset                (rst_controller_001_reset_out_reset),                                 //                   reset.reset
		.master_readdatavalid (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (pixel_buffer_dma_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (pixel_buffer_dma_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (pixel_buffer_dma_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (pixel_buffer_dma_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_dma_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_dma_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (pixel_buffer_dma_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (pixel_buffer_dma_avalon_pixel_source_data)                           //                        .data
	);

	Altera_UP_SD_Card_Avalon_Interface sd_card (
		.i_avalon_chip_select (mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (mm_interconnect_0_sd_card_avalon_sdcard_slave_address),     //                    .address
		.i_avalon_read        (mm_interconnect_0_sd_card_avalon_sdcard_slave_read),        //                    .read
		.i_avalon_write       (mm_interconnect_0_sd_card_avalon_sdcard_slave_write),       //                    .write
		.i_avalon_byteenable  (mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable),  //                    .byteenable
		.i_avalon_writedata   (mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata),   //                    .writedata
		.o_avalon_readdata    (mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata),    //                    .readdata
		.o_avalon_waitrequest (mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest), //                    .waitrequest
		.i_clock              (altpll_c0_clk),                                             //                 clk.clk
		.i_reset_n            (~rst_controller_001_reset_out_reset),                       //               reset.reset_n
		.b_SD_cmd             (sd_card_wire_b_SD_cmd),                                     //         conduit_end.export
		.b_SD_dat             (sd_card_wire_b_SD_dat),                                     //                    .export
		.b_SD_dat3            (sd_card_wire_b_SD_dat3),                                    //                    .export
		.o_SD_clock           (sd_card_wire_o_SD_clock)                                    //                    .export
	);

	Qsys_system_sdram sdram (
		.clk            (altpll_c0_clk),                            //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	Qsys_system_sysid sysid (
		.clock    (altpll_c0_clk),                                  //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	Qsys_system_timer timer (
		.clk        (altpll_c0_clk),                         //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	Qsys_system_vga_controller vga_controller (
		.clk           (altpll_c2_clk),                                           //                clk.clk
		.reset         (rst_controller_002_reset_out_reset),                      //              reset.reset
		.data          (dual_clock_buffer_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (dual_clock_buffer_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (dual_clock_buffer_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (dual_clock_buffer_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (dual_clock_buffer_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_controller_wire_CLK),                                 // external_interface.export
		.VGA_HS        (vga_controller_wire_HS),                                  //                   .export
		.VGA_VS        (vga_controller_wire_VS),                                  //                   .export
		.VGA_BLANK     (vga_controller_wire_BLANK),                               //                   .export
		.VGA_SYNC      (vga_controller_wire_SYNC),                                //                   .export
		.VGA_R         (vga_controller_wire_R),                                   //                   .export
		.VGA_G         (vga_controller_wire_G),                                   //                   .export
		.VGA_B         (vga_controller_wire_B)                                    //                   .export
	);

	Qsys_system_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (altpll_c0_clk),                                         //               clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                    //             reset.reset
		.stream_in_startofpacket  (pixel_buffer_dma_avalon_pixel_source_startofpacket),    //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_dma_avalon_pixel_source_endofpacket),      //                  .endofpacket
		.stream_in_valid          (pixel_buffer_dma_avalon_pixel_source_valid),            //                  .valid
		.stream_in_ready          (pixel_buffer_dma_avalon_pixel_source_ready),            //                  .ready
		.stream_in_data           (pixel_buffer_dma_avalon_pixel_source_data),             //                  .data
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)           //                  .data
	);

	Qsys_system_wifi_uart wifi_uart (
		.clk           (altpll_c0_clk),                                //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address       (mm_interconnect_0_wifi_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_wifi_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_wifi_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_wifi_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_wifi_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_wifi_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_wifi_uart_s1_readdata),      //                    .readdata
		.dataavailable (),                                             //                    .dataavailable
		.readyfordata  (),                                             //                    .readyfordata
		.rxd           (wifi_uart_wire_rxd),                           // external_connection.export
		.txd           (wifi_uart_wire_txd),                           //                    .export
		.cts_n         (wifi_uart_wire_cts_n),                         //                    .export
		.rts_n         (wifi_uart_wire_rts_n),                         //                    .export
		.irq           (irq_mapper_receiver2_irq)                      //                 irq.irq
	);

	Qsys_system_mm_interconnect_0 mm_interconnect_0 (
		.altpll_c0_clk                                            (altpll_c0_clk),                                                      //                                          altpll_c0.clk
		.clk_0_clk_clk                                            (clk_clk),                                                            //                                          clk_0_clk.clk
		.altpll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                     // altpll_inclk_interface_reset_reset_bridge_in_reset.reset
		.pixel_buffer_dma_reset_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),                                 //       pixel_buffer_dma_reset_reset_bridge_in_reset.reset
		.nios2_gen2_data_master_address                           (nios2_gen2_data_master_address),                                     //                             nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                       (nios2_gen2_data_master_waitrequest),                                 //                                                   .waitrequest
		.nios2_gen2_data_master_byteenable                        (nios2_gen2_data_master_byteenable),                                  //                                                   .byteenable
		.nios2_gen2_data_master_read                              (nios2_gen2_data_master_read),                                        //                                                   .read
		.nios2_gen2_data_master_readdata                          (nios2_gen2_data_master_readdata),                                    //                                                   .readdata
		.nios2_gen2_data_master_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                               //                                                   .readdatavalid
		.nios2_gen2_data_master_write                             (nios2_gen2_data_master_write),                                       //                                                   .write
		.nios2_gen2_data_master_writedata                         (nios2_gen2_data_master_writedata),                                   //                                                   .writedata
		.nios2_gen2_data_master_debugaccess                       (nios2_gen2_data_master_debugaccess),                                 //                                                   .debugaccess
		.nios2_gen2_instruction_master_address                    (nios2_gen2_instruction_master_address),                              //                      nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest                (nios2_gen2_instruction_master_waitrequest),                          //                                                   .waitrequest
		.nios2_gen2_instruction_master_read                       (nios2_gen2_instruction_master_read),                                 //                                                   .read
		.nios2_gen2_instruction_master_readdata                   (nios2_gen2_instruction_master_readdata),                             //                                                   .readdata
		.nios2_gen2_instruction_master_readdatavalid              (nios2_gen2_instruction_master_readdatavalid),                        //                                                   .readdatavalid
		.pixel_buffer_dma_avalon_pixel_dma_master_address         (pixel_buffer_dma_avalon_pixel_dma_master_address),                   //           pixel_buffer_dma_avalon_pixel_dma_master.address
		.pixel_buffer_dma_avalon_pixel_dma_master_waitrequest     (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),               //                                                   .waitrequest
		.pixel_buffer_dma_avalon_pixel_dma_master_read            (pixel_buffer_dma_avalon_pixel_dma_master_read),                      //                                                   .read
		.pixel_buffer_dma_avalon_pixel_dma_master_readdata        (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                  //                                                   .readdata
		.pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid   (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),             //                                                   .readdatavalid
		.pixel_buffer_dma_avalon_pixel_dma_master_lock            (pixel_buffer_dma_avalon_pixel_dma_master_lock),                      //                                                   .lock
		.altpll_pll_slave_address                                 (mm_interconnect_0_altpll_pll_slave_address),                         //                                   altpll_pll_slave.address
		.altpll_pll_slave_write                                   (mm_interconnect_0_altpll_pll_slave_write),                           //                                                   .write
		.altpll_pll_slave_read                                    (mm_interconnect_0_altpll_pll_slave_read),                            //                                                   .read
		.altpll_pll_slave_readdata                                (mm_interconnect_0_altpll_pll_slave_readdata),                        //                                                   .readdata
		.altpll_pll_slave_writedata                               (mm_interconnect_0_altpll_pll_slave_writedata),                       //                                                   .writedata
		.chaos_code_done_s1_address                               (mm_interconnect_0_chaos_code_done_s1_address),                       //                                 chaos_code_done_s1.address
		.chaos_code_done_s1_write                                 (mm_interconnect_0_chaos_code_done_s1_write),                         //                                                   .write
		.chaos_code_done_s1_readdata                              (mm_interconnect_0_chaos_code_done_s1_readdata),                      //                                                   .readdata
		.chaos_code_done_s1_writedata                             (mm_interconnect_0_chaos_code_done_s1_writedata),                     //                                                   .writedata
		.chaos_code_done_s1_chipselect                            (mm_interconnect_0_chaos_code_done_s1_chipselect),                    //                                                   .chipselect
		.chaos_code_reset_s1_address                              (mm_interconnect_0_chaos_code_reset_s1_address),                      //                                chaos_code_reset_s1.address
		.chaos_code_reset_s1_write                                (mm_interconnect_0_chaos_code_reset_s1_write),                        //                                                   .write
		.chaos_code_reset_s1_readdata                             (mm_interconnect_0_chaos_code_reset_s1_readdata),                     //                                                   .readdata
		.chaos_code_reset_s1_writedata                            (mm_interconnect_0_chaos_code_reset_s1_writedata),                    //                                                   .writedata
		.chaos_code_reset_s1_chipselect                           (mm_interconnect_0_chaos_code_reset_s1_chipselect),                   //                                                   .chipselect
		.chaos_code_shift_s1_address                              (mm_interconnect_0_chaos_code_shift_s1_address),                      //                                chaos_code_shift_s1.address
		.chaos_code_shift_s1_write                                (mm_interconnect_0_chaos_code_shift_s1_write),                        //                                                   .write
		.chaos_code_shift_s1_readdata                             (mm_interconnect_0_chaos_code_shift_s1_readdata),                     //                                                   .readdata
		.chaos_code_shift_s1_writedata                            (mm_interconnect_0_chaos_code_shift_s1_writedata),                    //                                                   .writedata
		.chaos_code_shift_s1_chipselect                           (mm_interconnect_0_chaos_code_shift_s1_chipselect),                   //                                                   .chipselect
		.chaos_code_step_s1_address                               (mm_interconnect_0_chaos_code_step_s1_address),                       //                                 chaos_code_step_s1.address
		.chaos_code_step_s1_write                                 (mm_interconnect_0_chaos_code_step_s1_write),                         //                                                   .write
		.chaos_code_step_s1_readdata                              (mm_interconnect_0_chaos_code_step_s1_readdata),                      //                                                   .readdata
		.chaos_code_step_s1_writedata                             (mm_interconnect_0_chaos_code_step_s1_writedata),                     //                                                   .writedata
		.chaos_code_step_s1_chipselect                            (mm_interconnect_0_chaos_code_step_s1_chipselect),                    //                                                   .chipselect
		.chaos_code_w_s1_address                                  (mm_interconnect_0_chaos_code_w_s1_address),                          //                                    chaos_code_w_s1.address
		.chaos_code_w_s1_write                                    (mm_interconnect_0_chaos_code_w_s1_write),                            //                                                   .write
		.chaos_code_w_s1_readdata                                 (mm_interconnect_0_chaos_code_w_s1_readdata),                         //                                                   .readdata
		.chaos_code_w_s1_writedata                                (mm_interconnect_0_chaos_code_w_s1_writedata),                        //                                                   .writedata
		.chaos_code_w_s1_chipselect                               (mm_interconnect_0_chaos_code_w_s1_chipselect),                       //                                                   .chipselect
		.chaos_code_x_s1_address                                  (mm_interconnect_0_chaos_code_x_s1_address),                          //                                    chaos_code_x_s1.address
		.chaos_code_x_s1_write                                    (mm_interconnect_0_chaos_code_x_s1_write),                            //                                                   .write
		.chaos_code_x_s1_readdata                                 (mm_interconnect_0_chaos_code_x_s1_readdata),                         //                                                   .readdata
		.chaos_code_x_s1_writedata                                (mm_interconnect_0_chaos_code_x_s1_writedata),                        //                                                   .writedata
		.chaos_code_x_s1_chipselect                               (mm_interconnect_0_chaos_code_x_s1_chipselect),                       //                                                   .chipselect
		.chaos_code_y_s1_address                                  (mm_interconnect_0_chaos_code_y_s1_address),                          //                                    chaos_code_y_s1.address
		.chaos_code_y_s1_write                                    (mm_interconnect_0_chaos_code_y_s1_write),                            //                                                   .write
		.chaos_code_y_s1_readdata                                 (mm_interconnect_0_chaos_code_y_s1_readdata),                         //                                                   .readdata
		.chaos_code_y_s1_writedata                                (mm_interconnect_0_chaos_code_y_s1_writedata),                        //                                                   .writedata
		.chaos_code_y_s1_chipselect                               (mm_interconnect_0_chaos_code_y_s1_chipselect),                       //                                                   .chipselect
		.chaos_code_z_s1_address                                  (mm_interconnect_0_chaos_code_z_s1_address),                          //                                    chaos_code_z_s1.address
		.chaos_code_z_s1_write                                    (mm_interconnect_0_chaos_code_z_s1_write),                            //                                                   .write
		.chaos_code_z_s1_readdata                                 (mm_interconnect_0_chaos_code_z_s1_readdata),                         //                                                   .readdata
		.chaos_code_z_s1_writedata                                (mm_interconnect_0_chaos_code_z_s1_writedata),                        //                                                   .writedata
		.chaos_code_z_s1_chipselect                               (mm_interconnect_0_chaos_code_z_s1_chipselect),                       //                                                   .chipselect
		.jtag_uart_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),              //                        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                //                                                   .write
		.jtag_uart_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                 //                                                   .read
		.jtag_uart_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),             //                                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),            //                                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),          //                                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),           //                                                   .chipselect
		.nios2_gen2_debug_mem_slave_address                       (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),               //                         nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                         (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),                 //                                                   .write
		.nios2_gen2_debug_mem_slave_read                          (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),                  //                                                   .read
		.nios2_gen2_debug_mem_slave_readdata                      (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),              //                                                   .readdata
		.nios2_gen2_debug_mem_slave_writedata                     (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),             //                                                   .writedata
		.nios2_gen2_debug_mem_slave_byteenable                    (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),            //                                                   .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest                   (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),           //                                                   .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess                   (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),           //                                                   .debugaccess
		.pio_key_s1_address                                       (mm_interconnect_0_pio_key_s1_address),                               //                                         pio_key_s1.address
		.pio_key_s1_write                                         (mm_interconnect_0_pio_key_s1_write),                                 //                                                   .write
		.pio_key_s1_readdata                                      (mm_interconnect_0_pio_key_s1_readdata),                              //                                                   .readdata
		.pio_key_s1_writedata                                     (mm_interconnect_0_pio_key_s1_writedata),                             //                                                   .writedata
		.pio_key_s1_chipselect                                    (mm_interconnect_0_pio_key_s1_chipselect),                            //                                                   .chipselect
		.pio_led_s1_address                                       (mm_interconnect_0_pio_led_s1_address),                               //                                         pio_led_s1.address
		.pio_led_s1_write                                         (mm_interconnect_0_pio_led_s1_write),                                 //                                                   .write
		.pio_led_s1_readdata                                      (mm_interconnect_0_pio_led_s1_readdata),                              //                                                   .readdata
		.pio_led_s1_writedata                                     (mm_interconnect_0_pio_led_s1_writedata),                             //                                                   .writedata
		.pio_led_s1_chipselect                                    (mm_interconnect_0_pio_led_s1_chipselect),                            //                                                   .chipselect
		.pio_wifi_reset_s1_address                                (mm_interconnect_0_pio_wifi_reset_s1_address),                        //                                  pio_wifi_reset_s1.address
		.pio_wifi_reset_s1_write                                  (mm_interconnect_0_pio_wifi_reset_s1_write),                          //                                                   .write
		.pio_wifi_reset_s1_readdata                               (mm_interconnect_0_pio_wifi_reset_s1_readdata),                       //                                                   .readdata
		.pio_wifi_reset_s1_writedata                              (mm_interconnect_0_pio_wifi_reset_s1_writedata),                      //                                                   .writedata
		.pio_wifi_reset_s1_chipselect                             (mm_interconnect_0_pio_wifi_reset_s1_chipselect),                     //                                                   .chipselect
		.pixel_buffer_avalon_sram_slave_address                   (mm_interconnect_0_pixel_buffer_avalon_sram_slave_address),           //                     pixel_buffer_avalon_sram_slave.address
		.pixel_buffer_avalon_sram_slave_write                     (mm_interconnect_0_pixel_buffer_avalon_sram_slave_write),             //                                                   .write
		.pixel_buffer_avalon_sram_slave_read                      (mm_interconnect_0_pixel_buffer_avalon_sram_slave_read),              //                                                   .read
		.pixel_buffer_avalon_sram_slave_readdata                  (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdata),          //                                                   .readdata
		.pixel_buffer_avalon_sram_slave_writedata                 (mm_interconnect_0_pixel_buffer_avalon_sram_slave_writedata),         //                                                   .writedata
		.pixel_buffer_avalon_sram_slave_byteenable                (mm_interconnect_0_pixel_buffer_avalon_sram_slave_byteenable),        //                                                   .byteenable
		.pixel_buffer_avalon_sram_slave_readdatavalid             (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdatavalid),     //                                                   .readdatavalid
		.pixel_buffer_dma_avalon_control_slave_address            (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address),    //              pixel_buffer_dma_avalon_control_slave.address
		.pixel_buffer_dma_avalon_control_slave_write              (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write),      //                                                   .write
		.pixel_buffer_dma_avalon_control_slave_read               (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read),       //                                                   .read
		.pixel_buffer_dma_avalon_control_slave_readdata           (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata),   //                                                   .readdata
		.pixel_buffer_dma_avalon_control_slave_writedata          (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata),  //                                                   .writedata
		.pixel_buffer_dma_avalon_control_slave_byteenable         (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable), //                                                   .byteenable
		.sd_card_avalon_sdcard_slave_address                      (mm_interconnect_0_sd_card_avalon_sdcard_slave_address),              //                        sd_card_avalon_sdcard_slave.address
		.sd_card_avalon_sdcard_slave_write                        (mm_interconnect_0_sd_card_avalon_sdcard_slave_write),                //                                                   .write
		.sd_card_avalon_sdcard_slave_read                         (mm_interconnect_0_sd_card_avalon_sdcard_slave_read),                 //                                                   .read
		.sd_card_avalon_sdcard_slave_readdata                     (mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata),             //                                                   .readdata
		.sd_card_avalon_sdcard_slave_writedata                    (mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata),            //                                                   .writedata
		.sd_card_avalon_sdcard_slave_byteenable                   (mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable),           //                                                   .byteenable
		.sd_card_avalon_sdcard_slave_waitrequest                  (mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest),          //                                                   .waitrequest
		.sd_card_avalon_sdcard_slave_chipselect                   (mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect),           //                                                   .chipselect
		.sdram_s1_address                                         (mm_interconnect_0_sdram_s1_address),                                 //                                           sdram_s1.address
		.sdram_s1_write                                           (mm_interconnect_0_sdram_s1_write),                                   //                                                   .write
		.sdram_s1_read                                            (mm_interconnect_0_sdram_s1_read),                                    //                                                   .read
		.sdram_s1_readdata                                        (mm_interconnect_0_sdram_s1_readdata),                                //                                                   .readdata
		.sdram_s1_writedata                                       (mm_interconnect_0_sdram_s1_writedata),                               //                                                   .writedata
		.sdram_s1_byteenable                                      (mm_interconnect_0_sdram_s1_byteenable),                              //                                                   .byteenable
		.sdram_s1_readdatavalid                                   (mm_interconnect_0_sdram_s1_readdatavalid),                           //                                                   .readdatavalid
		.sdram_s1_waitrequest                                     (mm_interconnect_0_sdram_s1_waitrequest),                             //                                                   .waitrequest
		.sdram_s1_chipselect                                      (mm_interconnect_0_sdram_s1_chipselect),                              //                                                   .chipselect
		.sysid_control_slave_address                              (mm_interconnect_0_sysid_control_slave_address),                      //                                sysid_control_slave.address
		.sysid_control_slave_readdata                             (mm_interconnect_0_sysid_control_slave_readdata),                     //                                                   .readdata
		.timer_s1_address                                         (mm_interconnect_0_timer_s1_address),                                 //                                           timer_s1.address
		.timer_s1_write                                           (mm_interconnect_0_timer_s1_write),                                   //                                                   .write
		.timer_s1_readdata                                        (mm_interconnect_0_timer_s1_readdata),                                //                                                   .readdata
		.timer_s1_writedata                                       (mm_interconnect_0_timer_s1_writedata),                               //                                                   .writedata
		.timer_s1_chipselect                                      (mm_interconnect_0_timer_s1_chipselect),                              //                                                   .chipselect
		.wifi_uart_s1_address                                     (mm_interconnect_0_wifi_uart_s1_address),                             //                                       wifi_uart_s1.address
		.wifi_uart_s1_write                                       (mm_interconnect_0_wifi_uart_s1_write),                               //                                                   .write
		.wifi_uart_s1_read                                        (mm_interconnect_0_wifi_uart_s1_read),                                //                                                   .read
		.wifi_uart_s1_readdata                                    (mm_interconnect_0_wifi_uart_s1_readdata),                            //                                                   .readdata
		.wifi_uart_s1_writedata                                   (mm_interconnect_0_wifi_uart_s1_writedata),                           //                                                   .writedata
		.wifi_uart_s1_begintransfer                               (mm_interconnect_0_wifi_uart_s1_begintransfer),                       //                                                   .begintransfer
		.wifi_uart_s1_chipselect                                  (mm_interconnect_0_wifi_uart_s1_chipselect)                           //                                                   .chipselect
	);

	Qsys_system_irq_mapper irq_mapper (
		.clk           (altpll_c0_clk),                      //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_gen2_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset),   // reset_in1.reset
		.clk            (altpll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_c2_clk),                        //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

endmodule
