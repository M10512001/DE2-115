	component Qsys_system is
		port (
			clk_clk                : in    std_logic                     := 'X';             -- clk
			pio_chaos_done_export  : in    std_logic                     := 'X';             -- export
			pio_chaos_reset_export : out   std_logic;                                        -- export
			pio_chaos_shift_export : out   std_logic_vector(31 downto 0);                    -- export
			pio_chaos_step_export  : out   std_logic;                                        -- export
			reset_reset_n          : in    std_logic                     := 'X';             -- reset_n
			sdram_clk_clk          : out   std_logic;                                        -- clk
			sdram_wire_addr        : out   std_logic_vector(12 downto 0);                    -- addr
			sdram_wire_ba          : out   std_logic_vector(1 downto 0);                     -- ba
			sdram_wire_cas_n       : out   std_logic;                                        -- cas_n
			sdram_wire_cke         : out   std_logic;                                        -- cke
			sdram_wire_cs_n        : out   std_logic;                                        -- cs_n
			sdram_wire_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- dq
			sdram_wire_dqm         : out   std_logic_vector(3 downto 0);                     -- dqm
			sdram_wire_ras_n       : out   std_logic;                                        -- ras_n
			sdram_wire_we_n        : out   std_logic;                                        -- we_n
			pio_chaos_x_export     : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			pio_chaos_y_export     : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			pio_chaos_z_export     : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			pio_chaos_w_export     : in    std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component Qsys_system;

	u0 : component Qsys_system
		port map (
			clk_clk                => CONNECTED_TO_clk_clk,                --             clk.clk
			pio_chaos_done_export  => CONNECTED_TO_pio_chaos_done_export,  --  pio_chaos_done.export
			pio_chaos_reset_export => CONNECTED_TO_pio_chaos_reset_export, -- pio_chaos_reset.export
			pio_chaos_shift_export => CONNECTED_TO_pio_chaos_shift_export, -- pio_chaos_shift.export
			pio_chaos_step_export  => CONNECTED_TO_pio_chaos_step_export,  --  pio_chaos_step.export
			reset_reset_n          => CONNECTED_TO_reset_reset_n,          --           reset.reset_n
			sdram_clk_clk          => CONNECTED_TO_sdram_clk_clk,          --       sdram_clk.clk
			sdram_wire_addr        => CONNECTED_TO_sdram_wire_addr,        --      sdram_wire.addr
			sdram_wire_ba          => CONNECTED_TO_sdram_wire_ba,          --                .ba
			sdram_wire_cas_n       => CONNECTED_TO_sdram_wire_cas_n,       --                .cas_n
			sdram_wire_cke         => CONNECTED_TO_sdram_wire_cke,         --                .cke
			sdram_wire_cs_n        => CONNECTED_TO_sdram_wire_cs_n,        --                .cs_n
			sdram_wire_dq          => CONNECTED_TO_sdram_wire_dq,          --                .dq
			sdram_wire_dqm         => CONNECTED_TO_sdram_wire_dqm,         --                .dqm
			sdram_wire_ras_n       => CONNECTED_TO_sdram_wire_ras_n,       --                .ras_n
			sdram_wire_we_n        => CONNECTED_TO_sdram_wire_we_n,        --                .we_n
			pio_chaos_x_export     => CONNECTED_TO_pio_chaos_x_export,     --     pio_chaos_x.export
			pio_chaos_y_export     => CONNECTED_TO_pio_chaos_y_export,     --     pio_chaos_y.export
			pio_chaos_z_export     => CONNECTED_TO_pio_chaos_z_export,     --     pio_chaos_z.export
			pio_chaos_w_export     => CONNECTED_TO_pio_chaos_w_export      --     pio_chaos_w.export
		);

